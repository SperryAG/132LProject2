----------------------------------------------------------------------------------
-- Create Date:    13:09:50 01/18/2016 
-- Module Name:    ALU_32Bit - Behavioral 
----------------------------------------------------------------------------------
----------------------------------------------------------------------------------
-- LIBRARIES / PACKAGES
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
----------------------------------------------------------------------------------
-- ENTITY
----------------------------------------------------------------------------------
ENTITY ALU_32Bit IS
	PORT( 
		Func_in    : IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
      A_in       : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
      B_in       : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
      O_out      : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		Branch_out : OUT STD_LOGIC;
		Jump_out   : OUT STD_LOGIC 
	);
END ALU_32Bit;
----------------------------------------------------------------------------------
-- ARCHITECTURE
----------------------------------------------------------------------------------
ARCHITECTURE Behavioral OF ALU_32Bit IS
BEGIN

END Behavioral;

